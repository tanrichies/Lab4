`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:26:45 03/02/2016 
// Design Name: 
// Module Name:    Led_Controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module led_controller(clk, reset, a7, a6, a5, a4, a3, a2 ,a1, seg_sel);
input 			clk, reset;
output 			a7, a6, a5, a4, a3, a2, a1, a0;
output 	[2:0]	seg_sel;
























endmodule
